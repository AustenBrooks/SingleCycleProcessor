----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/07/2021 07:12:52 PM
-- Design Name: 
-- Module Name: register_file - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity register_file is
    Port ( regSelReadA : in STD_LOGIC_VECTOR (4 downto 0);
           regSelReadB : in STD_LOGIC_VECTOR (4 downto 0);
           regSelWrite : in STD_LOGIC_VECTOR (4 downto 0);
           writeData : in STD_LOGIC_VECTOR (63 downto 0);
           regWrite : in STD_LOGIC;
           outA : out STD_LOGIC_VECTOR (63 downto 0);
           outB : out STD_LOGIC_VECTOR (63 downto 0));
end register_file;

architecture Behavioral of register_file is
type REG is array (0 to 31) of std_logic_vector(63 downto 0);
    signal registers : REG := (
    "0000000000000000000000000000000000000000000000000000000000000000", --X0
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000", --X10
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000", --X20
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000", --X30
    "0000000000000000000000000000000000000000000000000000000000000000");
begin
    process (regSelReadA, regSelReadB, regSelWrite, writeData, regWrite) is
        begin
        
        outA <= registers(to_integer(unsigned(regSelReadA)));
        outB <= registers(to_integer(unsigned(regSelReadB)));
        
        if regWrite = '1' then
            registers(to_integer(unsigned(regSelWrite))) <= writeData;
        end if;
    end process;
    

end Behavioral;
